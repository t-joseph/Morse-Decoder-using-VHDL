---------------------------------------------------------------------------------------
--------------------------Filename: mux.vhd - 12x1 MUX---------------------------------
---------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
---------------------------------------------------------------------------------------
ENTITY mux12x1 is
  PORT (data_i : IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
        sel_i  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	    y_o  : OUT STD_LOGIC);
  END mux12x1;
---------------------------------------------------------------------------------------

ARCHITECTURE a1 OF mux12x1 IS 

BEGIN 

  WITH sel_i SELECT
  y_o <= 
         '1' WHEN "0000",
         '0' WHEN "0001",     
         data_i(0) WHEN "0010",
         data_i(1) WHEN "0011",
         data_i(2) WHEN "0100",
         data_i(3) WHEN "0101",
         data_i(4) WHEN "0110",
         data_i(5) WHEN "0111",
         data_i(6) WHEN "1000", 
         data_i(7) WHEN "1001",
         '1' WHEN "1010",
         '1' WHEN "1011",
         '1' WHEN OTHERS;
END a1;
---------------------------------------------------------------------------------------