-----------------------------------------------------------------
---------------and2.vhd - 2 INPUT AND---------------------------
-----------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------------
ENTITY wgt_and2 IS
PORT (i1,i2:IN STD_LOGIC; o1:OUT STD_LOGIC);
END wgt_and2;
-----------------------------------------------------------------

ARCHITECTURE a1 OF wgt_and2 IS
BEGIN o1 <= i1 AND i2 AFTER 6 NS;
-----------------------------------------------------------------
END a1;
-----------------------------------------------------------------